module tb ();
    initial begin
        $dumpfile("dump.lxt");
        $dumpvars();
    end    
endmodule
